altclkctrl0_inst : altclkctrl0 PORT MAP (
		inclk	 => inclk_sig,
		outclk	 => outclk_sig
	);
