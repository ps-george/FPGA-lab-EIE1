lpm_counter5_inst : lpm_counter5 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
