bigcounter1_inst : bigcounter1 PORT MAP (
		aclr	 => aclr_sig,
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
